//I2C subordinate module. Work in progress.
