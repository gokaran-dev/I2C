//IC2 Subordinate modules 

